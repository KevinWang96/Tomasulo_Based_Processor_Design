/*
 * @Author: Yihao Wang
 * @Date: 2020-04-28 00:39:38
 * @LastEditTime: 2020-04-28 05:29:35
 * @LastEditors: Please set LastEditors
 * @Description: 
 *       a. Free Register List implemented using a sync FIFO
 *       b. Contact with DU: offering unused PID to DU during instruction dispatching
 *       c. Contact with CFC: also offering same unused PID to CFC during instruction dispatching
 *           and changing read pointer during flushing due miss branch prediction
 *       d. Contact with ROB: If an intruction graduated from ROB, it should return its old PID for Rd 
 *           back to FRL to ensure recycling of PID
 * @FilePath: /Tomasulo_3/Tomasulo_3_test1/projects/design/frl.v
 */
 `define FRL_DEPTH = 96 // 128 PIDs are needed but 32 of them are preinitialized in CFC (FRAT)
 `define FRL_WIDTH = 7 // since there are 128 locations in PRF (physical register file)
 module frl (
     clk, reset,
     dispatch_pid, pid_out,
     return_pid, pid_in,
     flush_frl, flush_frl_value
 );

    localparam FRL_PTR_WIDTH = `FRL_WIDTH + 1; // (n + 1)-bit pointer

    input dispatch_pid; // 1-bit dispath control signal and generated by DU
    output [0:`FRL_WIDTH - 1] pid_out; // PID dispatched from FRL
    output frl_empty; // no PID in frl, DU must stall dispatching

    input return_pid; // 1-bit return control signal and generated by ROB
    input [0:`FRL_WIDTH - 1] pid_in; // PID returned by ROB

    input flush_frl; // 1-bit flush control signal and generated by CFC
    input [0:FRL_PTR_WIDTH - 1] flush_frl_value; // flush value given by CFC

    // Instantiates a sync FIFO
    sync_fifo #(
        .DEPTH(`FRL_DEPTH),
        .WIDTH(`FRL_WIDTH),
        .PTR_WIDTH(FRL_PTR_WIDTH),
        .RESET_MODE(3) // using reset mode 3, reset FRL with PID #32 to PID #128
    )
    sync_fifo_inst
    (
        .clk(clk), .reset(reset),
        .r_en(dispatch_pid), .dout(pid_out), .empty(frl_empty),
        .w_en(return_pid), .din(pid_in), .full(),
        .w_fail(), .r_fail(),
        .change_r_ptr_en(flush_frl), .change_r_ptr_value(flush_frl_value),
        .change_w_ptr_en(1'b0), .change_w_ptr_value({FRL_PTR_WIDTH{1'b0}}) // don't need to flush write pointer
    );

 endmodule
 `undef FRL_WIDTH
 `undef FRL_DEPTH