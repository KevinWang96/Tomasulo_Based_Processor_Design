/*
 * @Author: Yihao Wang
 * @Date: 2020-05-01 01:43:21
 * @LastEditTime: 2020-05-01 06:18:12
 * @LastEditors: Please set LastEditors
 * @Description: 
 *      a. 32 X 41 Reorder Buffer which is a FIFO-based
 *      b. 41-bit ROB entry for register write instructions (ADD, ADDi, SUB, SLL, MULT, DIV, LW, JAL) :
 *          {cur_rd_PID(6-bit), pre_rd_PID(6-bit), rd_AID(5-bit), reg_wr(1-bit), mem_wr(1-bit), complete(1-bit), unused_field(21-bit)};
 *      c. 41-bit ROB entry for memory write instructions (SW) :
 *          {rs_PID(6-bit), sw_addr_part0(11-bit), reg_wr(1-bit), mem_wr(1-bit), complete(1-bit), sw_addr_part1(21-bit)};
 *      d. It has one write-only port, one random-access port and one read-only port;
 *          write-only port is used to form an ROB entry by DU;
 *          random-access port is used to change the information indexed by ROB tag given by CDB;
 *          read-only port is used by graduation logic to make an instruction graduate form ROB;
 * @FilePath: /Tomasulo_3_test1/projects/design/rob.v
 */
 `include "./design/params/rob_params.v" // include macro definition file
 module rob (
    clk, 
    reset,

    du_w_en,
    du_w_din,
    rob_full,
    rob_rob_tag,

    cdb_w_en,
    cdb_rob_tag, 
    cdb_reg_wr,
    cdb_w_sw_addr,
    cdb_mem_wr,

    cfc_flush,
    cfc_flush_rob_tag,

    gu_r_en,
    gu_r_dout,
    rob_empty
);

    input                               clk;                // positive triggering system
    input                               reset;              // sync reset

    input                               du_w_en;            // write enbale generated by DU
    input   [0:`ROB_WIDTH - 1]          du_w_din;           // write data in of DU
    output                              rob_full;           // full signal
    output  [0:`ROB_ROB_TAG_WIDTH - 1]  rob_rob_tag;        // ROB tag given to DU

    input                               cdb_w_en;           // write enable generated by CDB
    input   [0:`ROB_ROB_TAG_WIDTH - 1]  cdb_rob_tag;        // ROB tag used to index ROB
    input                               cdb_reg_wr;         // register write signal given by CDB
    input   [0:`ROB_SW_ADDR_WIDTH - 1]  cdb_w_sw_addr;      // SW address given by CDB
    input                               cdb_mem_wr;         // memory write signal given by CDB

    input                               cfc_flush;          // flush signal from CFC
    input   [0:`ROB_ROB_TAG_WIDTH - 1]  cfc_flush_rob_tag;  // flush ROB with rob_tag

    input                               gu_r_en;            // read enable generated by graduation unit
    output  [0:`ROB_WIDTH - 1]          gu_r_dout;          // read data out of graduation unit
    input                               rob_empty;          // emoty signal

    wire                                rob_full; 
    wire    [0:`ROB_ROB_TAG_WIDTH - 1]  rob_rob_tag;
    wire    [0:`ROB_WIDTH - 1]          gu_r_dout; 

    reg     [0:`ROB_PTR_WIDTH - 1]      w_ptr;              // write pointer
    reg     [0:`ROB_PTR_WIDTH - 1]      r_ptr;              // read pointer
    wire    [0:`ROB_PTR_WIDTH - 1]      diff;               // difference between w_ptr and r_ptr

    wire                                rob_w_en_q;         // qualified write enable
    wire                                rob_r_en_q;         // qualified read enable

    wire    [0:`ROB_PTR_WIDTH - 1]      rob_flush_value;    // the value need to be flushed into w_ptr

    reg     [0:`ROB_WIDTH - 1]          mem     [0:`ROB_DEPTH - 1]; // memory array

    assign  rob_w_en_q      =   (du_w_en && (!rob_full));       // generates qualified write enable 
    assign  rob_r_en_q      =   (gu_r_en && (!rob_empty));      // generates qualified read enable 
    
    assign  diff            =   w_ptr - r_ptr;                  // generates diff    
    assign  rob_full        =   (diff == `ROB_DEPTH);           // generates rob_full
    assign  rob_empty       =   (diff == 0);                    // generates rob_empty

    assign  rob_rob_tag     =   w_ptr[1:`ROB_PTR_WIDTH - 1];    // generates rob_rob_tag

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    assign  rob_flush_value =   (cfc_flush_rob_tag >= r_ptr[1:`ROB_PTR_WIDTH - 1]) ?           // ???????????????????????????
                                    {r_ptr[0], cfc_flush_rob_tag} :
                                    {~r_ptr[0], cfc_flush_rob_tag};                            // Not sure !!!!!!!!!!!! 
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

//// Data writing
    always @(posedge clk) begin
        if(reset) begin
            r_ptr <= `ROB_READ_PTR_INIT_VALUE;
            w_ptr <= `ROB_WRITE_PTR_INIT_VALUE;
        end
        else begin
            // We assume that it is impossible that DU and CDB access 
            // the same ROB location at the same clock

            if(cfc_flush) w_ptr <= rob_flush_value; // flush w_ptr has higher priority than writing
            else if(rob_w_en_q) begin
                mem[w_ptr[1:`ROB_PTR_WIDTH - 1]] <= du_w_din;
                w_ptr <= w_ptr + 1;
            end

            if(cdb_w_en) 
                case({cdb_reg_wr, cdb_mem_wr})
                    2'b00 : mem[cdb_rob_tag][`ROB_COMP_START_LOC] <= 1;
                    2'b01 : begin
                        mem[cdb_rob_tag][`ROB_SW_ADDR_PART0_START_LOC+:`ROB_SW_ADDR_PART0_WIDTH] 
                            <= cdb_w_sw_addr[0+:`ROB_SW_ADDR_PART0_WIDTH];
                        mem[cdb_rob_tag][`ROB_SW_ADDR_PART1_START_LOC+:`ROB_SW_ADDR_PART1_WIDTH] 
                            <= cdb_w_sw_addr[`ROB_SW_ADDR_PART0_WIDTH+:`ROB_SW_ADDR_PART1_WIDTH];
                        mem[cdb_rob_tag][`ROB_COMP_START_LOC] <= 1;
                    end
                    2'b10 : mem[cdb_rob_tag][`ROB_COMP_START_LOC] <= 1;
                    // default : // ilegal
                endcase

        end
    end

//// Data reading 
    always @(posedge clk) 
        if(rob_r_en_q) r_ptr <= r_ptr + 1;
    
    assign  gu_r_dout   =   (rob_r_en_q) ? mem[r_ptr[1:`ROB_PTR_WIDTH - 1]] : `ROB_READ_DATA_OUT_IDLE;
                        
 endmodule