/*
 * @Author: Yihao Wang
 * @Date: 2020-04-28 03:02:55
 * @LastEditTime: 2020-04-28 05:33:14
 * @LastEditors: Please set LastEditors
 * @Description: 
 *      a. 8 X 2 Branch prediction buffer using 2-bit predictor
 *      b. One read-only port used by DU to lookup
 *      c. One read-write port used by CDB to lookup and update
 * @FilePath: /Tomasulo_3/Tomasulo_3_test1/projects/design/bpb.v
 */
 `define DEPTH = 8
 `define WIDTH = 2
 module bpb #(
     parameter RESET_VALUE = 2'b10 // reset BPB with 2'10 (weakly taken)
 )
 (
     clk, reset, 
     du_branch, du_bpb_addr, bpb_branch_prediction_du,
     cdb_branch, cdb_branch_res, cdb_bpb_addr, bpb_branch_prediction_cdb
 );
    
    localparam BPB_ADDR = $clog2(`DEPTH);

    input clk, reset; // positive edge triggering and synchronous reset

    input du_branch; // 1-bit branch signal generated by Dispatching Unit
    input [0:BPB_ADDR - 1] du_bpb_addr; // used to index BPB by DU
    output reg bpb_branch_prediction_du; // 1-bit branch prediction used by DU

    input cdb_branch; // 1-bit branch signal generated by CDB
    input cdb_branch_res; // 1-bit branch results signal generated by CDB
                          // 1 means taken, 0 means not taken
    input [0:BPB_ADDR - 1] cdb_bpb_addr; // used to index BPB by CDB
    output reg bpb_branch_prediction_cdb; // 1-bit branch prediction used by CDB

    // Memory array 
    reg [0:`WIDTH - 1] mem [0:`DEPTH - 1];

//// Read-write port:
    // Reading 
    always @(*) // generates CDB brach prediction based on 2-bit predictor
    begin
        if(!cdb_branch) bpb_branch_prediction_cdb = 0;
        else
            case(mem[cdb_bpb_addr])
                2'b00 : bpb_branch_prediction_cdb = 0;
                2'b01 : bpb_branch_prediction_cdb = 0;
                2'b10 : bpb_branch_prediction_cdb = 1;
                2'b11 : bpb_branch_prediction_cdb = 1;
            endcase
    end
    // Writing
    reg [0:`WIDTH - 1] updated_predictor;
    always @(*) // generates the output of incrementer or decrementer used by saturate counter
    begin
        updated_predictor = mem[cdb_bpb_addr]; // if saturated, keep it as it is

        if( !( ((mem[cdb_bpb_addr] == 2'b11) && (cdb_branch_res)) 
            || ((mem[cdb_bpb_addr] == 2'b00) && (!cdb_branch_res)) ) // make sure counter is not saturate
        )
        begin
            if(cdb_branch_res) updated_predictor = mem[cdb_bpb_addr] + 1;
            else updated_predictor = mem[cdb_bpb_addr] - 1;
        end  
    end 

    always @(posedge clk) // update BPB using results of adder
    begin
        if(reset) 
        begin : reset_loop
            integer i;
            for(i = 0; i < `DEPTH; i = i + 1) mem[i] <= RESET_VALUE;
        end
        else
            if(cdb_branch) mem[cdb_bpb_addr] <= updated_predictor;
    end

//// Read-only port:
    wire [0:`WIDTH - 1] read_predictor; // supports internally forwarding
    assign read_predictor = (du_bpb_addr == cdb_bpb_addr) ? updated_predictor : mem[cdb_bpb_addr];

    always @(*) // generates DU brach prediction based on 2-bit predictor
    begin 
        if(!du_branch) bpb_branch_prediction_du = 0;
        else // if du_branch == 1
            case(read_predictor)
                2'b00 : bpb_branch_prediction_du = 0;
                2'b01 : bpb_branch_prediction_du = 0;
                2'b10 : bpb_branch_prediction_du = 1;
                2'b11 : bpb_branch_prediction_du = 1;
            endcase
    end

 endmodule
 `undef DEPTH
 `undef WIDTH